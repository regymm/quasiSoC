//`define SIMULATION

// clock freq
`define CLOCK_FREQ 62500000;
// CPU features
`define RV32M

// peripheral features
`define GPIO_EN
`define UART_EN
`define PSRAM_EN
`define SDCARD_EN
//`define CH375B_EN
`define VIDEO_EN
`define VIDEO_FALSEDIFFPAIR
`define IRQ_EN
//`define PS2_EN
//`define MMU_EN

`define SERIALBOOT_EN
`define UART_RST_EN
