//`define SIMULATION

//`define CLOCK_FREQ 50000000;

// peripheral features  
`define GPIO_EN
`define UART_EN
`define UART_RV_EN
`define SDRAM_EN
//`define BRAM_EN
//`define PSRAM_EN
//`define CACHE_EN
`define SDCARD_EN
//`define CH375B_EN
//`define VIDEO_EN
//`define IRQ_EN
//`define PS2_EN
//`define ETH_EN
//`define MMU_EN

//`define SERIALBOOT_EN
`define UART_RST_EN
