/**
 * File              : rv32a.v
 * License           : GPL-3.0-or-later
 * Author            : Peter Gu <github.com/regymm>
 * Date              : 2022.07.06
 * Last Modified Date: 2022.07.06
 */
`timescale 1ns / 1ps

module rv32a
	(
    );
endmodule
