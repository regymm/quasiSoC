//`define SIMULATION

// clock freq
`define CLOCK_FREQ 62500000;
// CPU features
`define RV32M
`define RV32A
`define IRQ_EN

// peripheral features
`define GPIO_EN
`define UART_EN
`define UART2_EN
`define PSRAM_EN
`define CACHE_EN
`define SDCARD_EN
//`define CH375B_EN
`define VIDEO_EN
`define VT100_EN
//`define LCD_EN
//`define PS2_EN
//`define ETH_EN
//`define MMU_EN

`define SERIALBOOT_EN
`define UART_RST_EN

//`define AXI_GPIO_TEST
